LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY rom IS
    PORT (
        clk : IN STD_LOGIC;
        address : IN unsigned (15 DOWNTO 0);
        data : OUT unsigned (15 DOWNTO 0)
    );
END rom;

ARCHITECTURE a_rom OF rom IS
    TYPE mem IS ARRAY (0 TO 255) OF unsigned (15 DOWNTO 0);
    CONSTANT content_rom : mem := (
        0 => B"0001_001_0_00100001",
        1 => B"0001_000_1_00000000",
        2 => B"0111_0000_000_1_0000",
        3 => B"0101_000_1_00000000",
        4 => B"1000_0000_001_0_0000",
        5 => B"1101_0000_11111101",
        6 => B"0001_000_1_00000010",
        7 => B"0001_010_0_00000010",
        8 => B"0011_0000_010_00000",
        9 => B"0010_011_0_000_1_0000",
        10 => B"0001_000_1_00000000",
        11 => B"0111_0000_011_0_0000",
        12 => B"0010_000_1_011_0_0000",
        13 => B"1000_0000_001_0_0000",
        14 => B"1011_0000_11111010",
        15 => B"0001_000_1_00000011",
        16 => B"0001_010_0_00000011",
        17 => B"0011_0000_010_00000",
        18 => B"0010_011_0_000_1_0000",
        19 => B"0001_000_1_00000000",
        20 => B"0111_0000_011_0_0000",
        21 => B"0010_000_1_011_0_0000",
        22 => B"1000_0000_001_0_0000",
        23 => B"1011_0000_11111010",
        24 => B"0001_000_1_00000101",
        25 => B"0001_010_0_00000101",
        26 => B"0011_0000_010_00000",
        27 => B"0010_011_0_000_1_0000",
        28 => B"0001_000_1_00000000",
        29 => B"0111_0000_011_0_0000",
        30 => B"0010_000_1_011_0_0000",
        31 => B"1000_0000_001_0_0000",
        32 => B"1011_0000_11111010",
        33 => B"0001_000_1_00000111",
        34 => B"0001_010_0_00000111",
        35 => B"0011_0000_010_00000",
        36 => B"0010_011_0_000_1_0000",
        37 => B"0001_000_1_00000000",
        38 => B"0111_0000_011_0_0000",
        39 => B"0010_000_1_011_0_0000",
        40 => B"1000_0000_001_0_0000",
        41 => B"1011_0000_11111010",
        42 => B"0001_000_1_00000010",
        43 => B"0110_110_0_000_1_0000",
        44 => B"0101_000_1_00000000",
        45 => B"1000_0000_001_0_0000",
        46 => B"1011_0000_11111101",
        
        OTHERS => (OTHERS => '0')
    );

BEGIN
    PROCESS (clk)
    BEGIN
        IF (rising_edge(clk)) THEN
            data <= content_rom(to_integer(address));
        END IF;
    END PROCESS;
END a_rom;